`timescale 1ns / 1ns

// registers are 32 bits in RV32
`define REG_SIZE 31

// RV opcodes are 7 bits
`define OPCODE_SIZE 6

module RegFile (
    input      [        4:0] rd,
    input      [`REG_SIZE:0] rd_data,
    input      [        4:0] rs1,
    output reg [`REG_SIZE:0] rs1_data,
    input      [        4:0] rs2,
    output reg [`REG_SIZE:0] rs2_data,
    input                    clk,
    input                    we,
    input                    rst
);
    localparam NumRegs = 32;
    reg [`REG_SIZE:0] regs[0:NumRegs-1];
    integer i;

    // --- Asynchronous Read ---
    // x0 is always hardwired to 0
    always @(*) begin
        rs1_data = (rs1 == 5'd0) ? 32'd0 : regs[rs1];
        rs2_data = (rs2 == 5'd0) ? 32'd0 : regs[rs2];
    end

    // --- Synchronous Write ---
    always @(posedge clk) begin
        if (rst) begin
            for (i = 0; i < NumRegs; i = i + 1) begin
                regs[i] <= 32'd0;
            end
        end else if (we && (rd != 5'd0)) begin
            regs[rd] <= rd_data;
        end
    end

endmodule

module DatapathSingleCycle (
    input                    clk,
    input                    rst,
    output reg               halt,
    output     [`REG_SIZE:0] pc_to_imem,
    input      [`REG_SIZE:0] inst_from_imem,
    // addr_to_dmem is a read-write port
    output reg [`REG_SIZE:0] addr_to_dmem,
    input      [`REG_SIZE:0] load_data_from_dmem,
    output reg [`REG_SIZE:0] store_data_to_dmem,
    output reg [        3:0] store_we_to_dmem
);
    // components of the instruction
    wire [           6:0] inst_funct7;
    wire [           4:0] inst_rs2;
    wire [           4:0] inst_rs1;
    wire [           2:0] inst_funct3;
    wire [           4:0] inst_rd;
    wire [`OPCODE_SIZE:0] inst_opcode;

    // split R-type instruction - see section 2.2 of RiscV spec
    assign {inst_funct7, inst_rs2, inst_rs1, inst_funct3, inst_rd, inst_opcode} = inst_from_imem;

    // setup for I, S, B & J type instructions
    // I - short immediates and loads
    wire [11:0] imm_i;
    assign imm_i = inst_from_imem[31:20];
    wire [ 4:0] imm_shamt = inst_from_imem[24:20];

    // S - stores
    wire [11:0] imm_s;
    assign imm_s = {inst_funct7, inst_rd};

    // B - conditionals
    wire [12:0] imm_b;
    assign {imm_b[12], imm_b[10:1], imm_b[11], imm_b[0]} = {inst_funct7, inst_rd, 1'b0};

    // J - unconditional jumps
    wire [20:0] imm_j;
    assign {imm_j[20], imm_j[10:1], imm_j[11], imm_j[19:12], imm_j[0]} = {inst_from_imem[31:12], 1'b0};

    // U - Upper immediate (LUI, AUIPC) - Missing from skeleton, added here
    wire [31:0] imm_u;
    assign imm_u = {inst_from_imem[31:12], 12'b0};

    wire [`REG_SIZE:0] imm_i_sext = {{20{imm_i[11]}}, imm_i[11:0]};
    wire [`REG_SIZE:0] imm_s_sext = {{20{imm_s[11]}}, imm_s[11:0]};
    wire [`REG_SIZE:0] imm_b_sext = {{19{imm_b[12]}}, imm_b[12:0]};
    wire [`REG_SIZE:0] imm_j_sext = {{11{imm_j[20]}}, imm_j[20:0]};

    // opcodes - see section 19 of RiscV spec
    localparam [`OPCODE_SIZE:0] OpLoad    = 7'b00_000_11;
    localparam [`OPCODE_SIZE:0] OpStore   = 7'b01_000_11;
    localparam [`OPCODE_SIZE:0] OpBranch  = 7'b11_000_11;
    localparam [`OPCODE_SIZE:0] OpJalr    = 7'b11_001_11;
    localparam [`OPCODE_SIZE:0] OpMiscMem = 7'b00_011_11;
    localparam [`OPCODE_SIZE:0] OpJal     = 7'b11_011_11;
    localparam [`OPCODE_SIZE:0] OpRegImm  = 7'b00_100_11;
    localparam [`OPCODE_SIZE:0] OpRegReg  = 7'b01_100_11;
    localparam [`OPCODE_SIZE:0] OpEnviron = 7'b11_100_11;
    localparam [`OPCODE_SIZE:0] OpAuipc   = 7'b00_101_11;
    localparam [`OPCODE_SIZE:0] OpLui     = 7'b01_101_11;

    wire inst_lui    = (inst_opcode == OpLui    );
    wire inst_auipc  = (inst_opcode == OpAuipc  );
    wire inst_jal    = (inst_opcode == OpJal    );
    wire inst_jalr   = (inst_opcode == OpJalr   );
    wire inst_beq    = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b000);
    wire inst_bne    = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b001);
    wire inst_blt    = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b100);
    wire inst_bge    = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b101);
    wire inst_bltu   = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b110);
    wire inst_bgeu   = (inst_opcode == OpBranch ) & (inst_from_imem[14:12] == 3'b111);
    wire inst_lb     = (inst_opcode == OpLoad   ) & (inst_from_imem[14:12] == 3'b000);
    wire inst_lh     = (inst_opcode == OpLoad   ) & (inst_from_imem[14:12] == 3'b001);
    wire inst_lw     = (inst_opcode == OpLoad   ) & (inst_from_imem[14:12] == 3'b010);
    wire inst_lbu    = (inst_opcode == OpLoad   ) & (inst_from_imem[14:12] == 3'b100);
    wire inst_lhu    = (inst_opcode == OpLoad   ) & (inst_from_imem[14:12] == 3'b101);
    wire inst_sb     = (inst_opcode == OpStore  ) & (inst_from_imem[14:12] == 3'b000);
    wire inst_sh     = (inst_opcode == OpStore  ) & (inst_from_imem[14:12] == 3'b001);
    wire inst_sw     = (inst_opcode == OpStore  ) & (inst_from_imem[14:12] == 3'b010);
    wire inst_addi   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b000);
    wire inst_slti   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b010);
    wire inst_sltiu  = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b011);
    wire inst_xori   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b100);
    wire inst_ori    = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b110);
    wire inst_andi   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b111);
    wire inst_slli   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b001) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_srli   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b101) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_srai   = (inst_opcode == OpRegImm ) & (inst_from_imem[14:12] == 3'b101) & (inst_from_imem[31:25] == 7'b0100000);
    wire inst_add    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b000) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_sub    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b000) & (inst_from_imem[31:25] == 7'b0100000);
    wire inst_sll    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b001) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_slt    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b010) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_sltu   = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b011) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_xor    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b100) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_srl    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b101) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_sra    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b101) & (inst_from_imem[31:25] == 7'b0100000);
    wire inst_or     = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b110) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_and    = (inst_opcode == OpRegReg ) & (inst_from_imem[14:12] == 3'b111) & (inst_from_imem[31:25] == 7'd0      );
    wire inst_mul    = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b000    );
    wire inst_mulh   = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b001    );
    wire inst_mulhsu = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b010    );
    wire inst_mulhu  = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b011    );
    wire inst_div    = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b100    );
    wire inst_divu   = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b101    );
    wire inst_rem    = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b110    );
    wire inst_remu   = (inst_opcode == OpRegReg ) & (inst_from_imem[31:25] == 7'd1  ) & (inst_from_imem[14:12] == 3'b111    );
    wire inst_ecall  = (inst_opcode == OpEnviron) & (inst_from_imem[31:7] == 25'd0  );
    wire inst_fence  = (inst_opcode == OpMiscMem);

    // program counter
    reg [`REG_SIZE:0] pcNext, pcCurrent;
    always @(posedge clk) begin
        if (rst) begin
            pcCurrent <= 32'd0;
        end else begin
            pcCurrent <= pcNext;
        end
    end
    assign pc_to_imem = pcCurrent;

    // cycle/inst counters
    reg [`REG_SIZE:0] cycles_current, num_inst_current;
    always @(posedge clk) begin
        if (rst) begin
            cycles_current <= 0;
            num_inst_current <= 0;
        end else begin
            cycles_current <= cycles_current + 1;
            if (!rst) begin
                num_inst_current <= num_inst_current + 1;
            end
        end
    end

    // --- REGISTER FILE ---
    wire [`REG_SIZE:0] rs1_data;
    wire [`REG_SIZE:0] rs2_data;
    reg [`REG_SIZE:0] rd_data_mux; // Data to write to RD
    reg rf_we_mux;                 // Write Enable mux

    RegFile rf (
        .clk      (clk),
        .rst      (rst),
        .we       (rf_we_mux),
        .rd       (inst_rd),
        .rd_data  (rd_data_mux),
        .rs1      (inst_rs1),
        .rs2      (inst_rs2),
        .rs1_data (rs1_data),
        .rs2_data (rs2_data)
    );

    // --- CLA ADDER ---
    wire [31:0] cla_op_a;
    wire [31:0] cla_op_b;
    wire [31:0] cla_sum;
    wire cla_sub_ctrl; // 1 for subtraction (invert B + cin)

    // For SUB, we invert B and add 1 (Cin). For ADD, we keep B and Cin=0.
    assign cla_op_a = rs1_data;
    // B operand is RS2 for R-type, Immediate for I-type
    assign cla_op_b = (inst_opcode == OpRegReg) ? rs2_data : imm_i_sext;
    // Control subtraction (only used for SUB instruction here, branch comparison is separate for simplicity)
    assign cla_sub_ctrl = inst_sub;

    cla my_cla (
        .a   (cla_op_a),
        .b   (cla_sub_ctrl ? ~cla_op_b : cla_op_b),
        .cin (cla_sub_ctrl),
        .sum (cla_sum)
    );

    // --- DIVIDER ---
    wire [31:0] div_rem_out;
    wire [31:0] div_quot_out;
    divider_unsigned my_div (
        .i_dividend (rs1_data),
        .i_divisor  (rs2_data),
        .o_remainder(div_rem_out),
        .o_quotient (div_quot_out)
    );

    // --- Control Logic & Datapath Muxes ---
    reg illegal_inst;

    always @(*) begin
        // Defaults to prevent latches
        illegal_inst = 1'b0;
        halt = 1'b0;
        pcNext = pcCurrent + 32'd4;
        rf_we_mux = 1'b0;
        rd_data_mux = 32'd0;
        addr_to_dmem = 32'd0;
        store_data_to_dmem = 32'd0;
        store_we_to_dmem = 4'b0000;

        case (inst_opcode)
            OpLui: begin
                rf_we_mux = 1'b1;
                rd_data_mux = imm_u;
            end
            OpAuipc: begin
                rf_we_mux = 1'b1;
                rd_data_mux = pcCurrent + imm_u; // Can use + operator per specs
            end
            OpJal: begin
                rf_we_mux = 1'b1;
                rd_data_mux = pcCurrent + 32'd4;
                pcNext = pcCurrent + imm_j_sext;
            end
            OpJalr: begin
                rf_we_mux = 1'b1;
                rd_data_mux = pcCurrent + 32'd4;
                // JALR target: (rs1 + offset) & ~1
                pcNext = (rs1_data + imm_i_sext) & ~32'd1;
            end
            OpBranch: begin
                // Branch Logic
                // Note: Comparisons done behaviorally for simplicity/timing
                if (inst_beq && (rs1_data == rs2_data)) pcNext = pcCurrent + imm_b_sext;
                else if (inst_bne && (rs1_data != rs2_data)) pcNext = pcCurrent + imm_b_sext;
                else if (inst_blt && ($signed(rs1_data) < $signed(rs2_data))) pcNext = pcCurrent + imm_b_sext;
                else if (inst_bge && ($signed(rs1_data) >= $signed(rs2_data))) pcNext = pcCurrent + imm_b_sext;
                else if (inst_bltu && (rs1_data < rs2_data)) pcNext = pcCurrent + imm_b_sext;
                else if (inst_bgeu && (rs1_data >= rs2_data)) pcNext = pcCurrent + imm_b_sext;
            end
            OpLoad: begin
                addr_to_dmem = rs1_data + imm_i_sext;
                rf_we_mux = 1'b1;
                // Handling sub-word loads
                case (inst_from_imem[14:12]) // funct3
                    3'b000: begin // LB
                        case(addr_to_dmem[1:0])
                           2'b00: rd_data_mux = {{24{load_data_from_dmem[7]}}, load_data_from_dmem[7:0]};
                           2'b01: rd_data_mux = {{24{load_data_from_dmem[15]}}, load_data_from_dmem[15:8]};
                           2'b10: rd_data_mux = {{24{load_data_from_dmem[23]}}, load_data_from_dmem[23:16]};
                           2'b11: rd_data_mux = {{24{load_data_from_dmem[31]}}, load_data_from_dmem[31:24]};
                        endcase
                    end
                    3'b001: begin // LH
                        case(addr_to_dmem[1:0])
                           2'b00: rd_data_mux = {{16{load_data_from_dmem[15]}}, load_data_from_dmem[15:0]};
                           2'b10: rd_data_mux = {{16{load_data_from_dmem[31]}}, load_data_from_dmem[31:16]};
                           default: rd_data_mux = 32'd0; // Unaligned
                        endcase
                    end
                    3'b010: rd_data_mux = load_data_from_dmem; // LW
                    3'b100: begin // LBU
                        case(addr_to_dmem[1:0])
                           2'b00: rd_data_mux = {24'd0, load_data_from_dmem[7:0]};
                           2'b01: rd_data_mux = {24'd0, load_data_from_dmem[15:8]};
                           2'b10: rd_data_mux = {24'd0, load_data_from_dmem[23:16]};
                           2'b11: rd_data_mux = {24'd0, load_data_from_dmem[31:24]};
                        endcase
                    end
                    3'b101: begin // LHU
                        case(addr_to_dmem[1:0])
                           2'b00: rd_data_mux = {16'd0, load_data_from_dmem[15:0]};
                           2'b10: rd_data_mux = {16'd0, load_data_from_dmem[31:16]};
                           default: rd_data_mux = 32'd0; // Unaligned
                        endcase
                    end
                    default: rd_data_mux = load_data_from_dmem;
                endcase
            end
            OpStore: begin
                addr_to_dmem = rs1_data + imm_s_sext;
                store_data_to_dmem = rs2_data << (8 * addr_to_dmem[1:0]); // Shift data to correct byte pos
                // Write Enable Logic based on funct3 and address alignment
                if (inst_sb)      store_we_to_dmem = 4'b0001 << addr_to_dmem[1:0];
                else if (inst_sh) store_we_to_dmem = 4'b0011 << addr_to_dmem[1:0];
                else if (inst_sw) store_we_to_dmem = 4'b1111;
            end
            OpRegImm: begin
                rf_we_mux = 1'b1;
                // ADDI uses CLA
                if (inst_addi) rd_data_mux = cla_sum;
                // Others use behavioural operators
                else if (inst_slti) rd_data_mux = ($signed(rs1_data) < $signed(imm_i_sext)) ? 32'd1 : 32'd0;
                else if (inst_sltiu) rd_data_mux = (rs1_data < imm_i_sext) ? 32'd1 : 32'd0;
                else if (inst_xori) rd_data_mux = rs1_data ^ imm_i_sext;
                else if (inst_ori)  rd_data_mux = rs1_data | imm_i_sext;
                else if (inst_andi) rd_data_mux = rs1_data & imm_i_sext;
                else if (inst_slli) rd_data_mux = rs1_data << imm_shamt;
                else if (inst_srli) rd_data_mux = rs1_data >> imm_shamt;
                else if (inst_srai) rd_data_mux = $signed(rs1_data) >>> imm_shamt;
            end
            OpRegReg: begin
                rf_we_mux = 1'b1;
                // ADD/SUB use CLA
                if (inst_add || inst_sub) rd_data_mux = cla_sum;
                // DIV/REM use Divider
                else if (inst_div)  rd_data_mux = ($signed(rs1_data) == -2147483648 && $signed(rs2_data) == -1) ? -2147483648 : 
                                                  (rs2_data == 0) ? -1 : ($signed(rs1_data) / $signed(rs2_data)); // Signed Div logic
                else if (inst_divu) rd_data_mux = div_quot_out; // Unsigned (Using your module)
                else if (inst_rem)  rd_data_mux = ($signed(rs1_data) == -2147483648 && $signed(rs2_data) == -1) ? 0 : 
                                                  (rs2_data == 0) ? rs1_data : ($signed(rs1_data) % $signed(rs2_data));
                else if (inst_remu) rd_data_mux = div_rem_out;  // Unsigned (Using your module)
                // Logical / Shift / Mul
                else if (inst_sll)  rd_data_mux = rs1_data << rs2_data[4:0];
                else if (inst_slt)  rd_data_mux = ($signed(rs1_data) < $signed(rs2_data)) ? 32'd1 : 32'd0;
                else if (inst_sltu) rd_data_mux = (rs1_data < rs2_data) ? 32'd1 : 32'd0;
                else if (inst_xor)  rd_data_mux = rs1_data ^ rs2_data;
                else if (inst_srl)  rd_data_mux = rs1_data >> rs2_data[4:0];
                else if (inst_sra)  rd_data_mux = $signed(rs1_data) >>> rs2_data[4:0];
                else if (inst_or)   rd_data_mux = rs1_data | rs2_data;
                else if (inst_and)  rd_data_mux = rs1_data & rs2_data;
                else if (inst_mul)  rd_data_mux = rs1_data * rs2_data;
                else if (inst_mulh)   rd_data_mux = 32'(($signed({{32{rs1_data[31]}}, rs1_data}) * $signed({{32{rs2_data[31]}}, rs2_data})) >> 32);
		else if (inst_mulhsu) rd_data_mux = 32'(($signed({{32{rs1_data[31]}}, rs1_data}) * $signed({32'd0, rs2_data})) >> 32);
		else if (inst_mulhu)  rd_data_mux = 32'(({{32'd0}, rs1_data} * {{32'd0}, rs2_data}) >> 32);
            end
            OpEnviron: begin
                if (inst_ecall) halt = 1'b1;
            end
            OpMiscMem: begin
                // FENCE - No op for this lab
            end
            default: begin
                illegal_inst = 1'b1;
            end
        endcase
    end

endmodule

/* A memory module that supports 1-cycle reads and writes */
module MemorySingleCycle #(
    parameter NUM_WORDS = 8192
) (
    input                    rst,
    input                    clock_mem,
    input      [`REG_SIZE:0] pc_to_imem,
    output reg [`REG_SIZE:0] inst_from_imem,
    input      [`REG_SIZE:0] addr_to_dmem,
    output reg [`REG_SIZE:0] load_data_from_dmem,
    input      [`REG_SIZE:0] store_data_to_dmem,
    input      [        3:0] store_we_to_dmem
);
    reg [`REG_SIZE:0] mem_array[0:NUM_WORDS-1];

    initial begin
        $readmemh("mem_initial_contents.hex", mem_array);
    end

    localparam AddrMsb = $clog2(NUM_WORDS) + 1;
    localparam AddrLsb = 2;

    always @(posedge clock_mem) begin
        inst_from_imem <= mem_array[{pc_to_imem[AddrMsb:AddrLsb]}];
    end

    always @(negedge clock_mem) begin
        if (store_we_to_dmem[0]) mem_array[addr_to_dmem[AddrMsb:AddrLsb]][7:0]   <= store_data_to_dmem[7:0];
        if (store_we_to_dmem[1]) mem_array[addr_to_dmem[AddrMsb:AddrLsb]][15:8]  <= store_data_to_dmem[15:8];
        if (store_we_to_dmem[2]) mem_array[addr_to_dmem[AddrMsb:AddrLsb]][23:16] <= store_data_to_dmem[23:16];
        if (store_we_to_dmem[3]) mem_array[addr_to_dmem[AddrMsb:AddrLsb]][31:24] <= store_data_to_dmem[31:24];

        load_data_from_dmem <= mem_array[{addr_to_dmem[AddrMsb:AddrLsb]}];
    end
endmodule

module Processor (
    input  clock_proc,
    input  clock_mem,
    input  rst,
    output halt
);
    wire [`REG_SIZE:0] pc_to_imem, inst_from_imem, mem_data_addr, mem_data_loaded_value, mem_data_to_write;
    wire [        3:0] mem_data_we;
    wire [(8*32)-1:0] test_case;

    MemorySingleCycle #(
        .NUM_WORDS(8192)
    ) memory (
        .rst                 (rst),
        .clock_mem           (clock_mem),
        .pc_to_imem          (pc_to_imem),
        .inst_from_imem      (inst_from_imem),
        .addr_to_dmem        (mem_data_addr),
        .load_data_from_dmem (mem_data_loaded_value),
        .store_data_to_dmem  (mem_data_to_write),
        .store_we_to_dmem    (mem_data_we)
    );

    DatapathSingleCycle datapath (
        .clk                 (clock_proc),
        .rst                 (rst),
        .pc_to_imem          (pc_to_imem),
        .inst_from_imem      (inst_from_imem),
        .addr_to_dmem        (mem_data_addr),
        .store_data_to_dmem  (mem_data_to_write),
        .store_we_to_dmem    (mem_data_we),
        .load_data_from_dmem (mem_data_loaded_value),
        .halt                (halt)
    );
endmodule
